module top_level_controller(
    input IN1,IN2,IN3,IN4,
    ENA,ENB,
    input [6:0] seg,
    input [3:0] an
);



endmodule
